VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO  tt_um_isshuwakita_r2r_dac
  CLASS BLOCK ;
  FOREIGN  tt_um_isshuwakita_r2r_dac ;
  ORIGIN -1.000 -5.000 ;
  SIZE 5.000 BY 215.760 ;
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
END  tt_um_isshuwakita_r2r_dac
END LIBRARY

