magic
tech sky130A
magscale 1 2
timestamp 1724825786
<< viali >>
rect 19426 738 19660 994
rect 19656 200 19738 352
rect 19172 -36 19386 184
rect 23030 28 23242 244
rect 26998 30 27194 266
rect 27970 246 28046 354
rect 30338 256 30524 470
rect 14912 -336 15180 -54
rect 28208 -1998 28442 -1636
<< metal1 >>
rect 19420 994 19666 1006
rect 19416 738 19426 994
rect 19660 738 19670 994
rect 19420 726 19666 738
rect 19486 600 19610 726
rect 19486 504 19618 600
rect 20080 584 20164 594
rect 19488 364 19618 504
rect 20068 572 23816 584
rect 27590 578 27774 584
rect 23968 574 27774 578
rect 23968 572 30754 574
rect 20068 504 30754 572
rect 20068 470 27774 504
rect 20068 454 24222 470
rect 19488 352 19744 364
rect 19488 200 19656 352
rect 19738 200 19744 352
rect 20080 342 20164 454
rect 23698 408 24222 454
rect 19822 336 20226 342
rect 19822 234 20332 336
rect 23698 334 24266 408
rect 27572 398 27774 470
rect 30244 470 30698 504
rect 27572 386 27918 398
rect 23698 320 24176 334
rect 27396 332 27918 386
rect 27964 358 28052 366
rect 27964 354 28484 358
rect 27396 326 27894 332
rect 23024 244 23248 256
rect 19498 196 19744 200
rect 19166 184 19392 196
rect 19650 188 19744 196
rect 19162 -36 19172 184
rect 19386 114 19396 184
rect 19894 138 20074 234
rect 20152 226 20332 234
rect 19386 56 19852 114
rect 19386 -36 19396 56
rect 20112 54 20168 112
rect 14906 -54 15186 -42
rect 19166 -48 19392 -36
rect 19898 -54 20078 34
rect 23020 28 23030 244
rect 23242 206 23252 244
rect 23838 230 24018 320
rect 27396 314 27818 326
rect 26992 266 27200 278
rect 23242 152 23786 206
rect 24048 152 24108 210
rect 23242 28 23252 152
rect 23836 42 24016 136
rect 23782 38 24112 42
rect 23024 16 23248 28
rect 23638 -22 24212 38
rect 26988 30 26998 266
rect 27194 204 27204 266
rect 27632 228 27818 314
rect 27964 246 27970 354
rect 28046 246 28484 354
rect 30244 348 30338 470
rect 27964 244 28484 246
rect 30288 256 30338 348
rect 30524 348 30698 470
rect 30524 256 30628 348
rect 27964 234 28052 244
rect 27194 140 27600 204
rect 27864 146 27924 208
rect 27194 30 27204 140
rect 27642 38 27822 130
rect 26992 18 27200 30
rect 27440 -22 28014 38
rect 14902 -336 14912 -54
rect 15180 -226 15190 -54
rect 19704 -114 20278 -54
rect 15180 -336 15200 -226
rect 14906 -348 15200 -336
rect 14914 -376 15200 -348
rect 19854 -376 20108 -114
rect 14914 -392 20108 -376
rect 23790 -392 24086 -22
rect 14914 -404 24086 -392
rect 27604 -404 27894 -22
rect 14914 -532 27894 -404
rect 14914 -562 20108 -532
rect 23786 -540 27894 -532
rect 27604 -550 27894 -540
rect 14914 -566 15200 -562
rect 19854 -568 20108 -562
rect 28236 -742 28452 244
rect 30288 200 30628 256
rect 28222 -1086 28452 -742
rect 28222 -1624 28448 -1086
rect 28202 -1636 28448 -1624
rect 28198 -1998 28208 -1636
rect 28442 -1998 28452 -1636
rect 28202 -2010 28448 -1998
<< via1 >>
rect 19426 738 19660 994
rect 19172 -36 19386 184
rect 23030 28 23242 244
rect 26998 30 27194 266
rect 30338 256 30524 470
rect 14912 -336 15180 -54
rect 28208 -1998 28442 -1636
<< metal2 >>
rect 19426 994 19660 1004
rect 19426 728 19660 738
rect 30338 470 30524 480
rect 26998 266 27194 276
rect 23030 244 23242 254
rect 19172 184 19386 194
rect 23030 18 23242 28
rect 30338 246 30524 256
rect 26998 20 27194 30
rect 14912 -54 15180 -44
rect 19172 -46 19386 -36
rect 14912 -346 15180 -336
rect 28208 -1636 28442 -1626
rect 28208 -2008 28442 -1998
<< via2 >>
rect 19426 738 19660 994
rect 19172 -36 19386 184
rect 23030 28 23242 244
rect 26998 30 27194 266
rect 30338 256 30524 470
rect 14912 -336 15180 -54
rect 28208 -1998 28442 -1636
<< metal3 >>
rect 19416 994 19670 999
rect 19416 738 19426 994
rect 19660 738 19670 994
rect 19416 733 19670 738
rect 30328 470 30534 475
rect 23020 244 23252 249
rect 19162 184 19396 189
rect 19162 -36 19172 184
rect 19386 -36 19396 184
rect 23020 28 23030 244
rect 23242 28 23252 244
rect 23020 23 23252 28
rect 26974 20 26984 276
rect 27214 20 27224 276
rect 30328 256 30338 470
rect 30524 256 30534 470
rect 30328 251 30534 256
rect 19162 -41 19396 -36
rect 14902 -54 15190 -49
rect 14902 -336 14912 -54
rect 15180 -336 15190 -54
rect 14902 -341 15190 -336
rect 28198 -1636 28452 -1631
rect 28198 -1998 28208 -1636
rect 28442 -1998 28452 -1636
rect 28198 -2003 28452 -1998
<< via3 >>
rect 19426 738 19660 994
rect 19172 -36 19386 184
rect 23030 28 23242 244
rect 26984 266 27214 276
rect 26984 30 26998 266
rect 26998 30 27194 266
rect 27194 30 27214 266
rect 26984 20 27214 30
rect 30338 256 30524 470
rect 14912 -336 15180 -54
rect 28208 -1998 28442 -1636
<< metal4 >>
rect 200 1712 600 44152
rect 800 2044 1200 44152
rect 198 1000 600 1712
rect 732 1250 19616 2044
rect 732 1160 19618 1250
rect 800 1000 1200 1160
rect 19248 1014 19618 1160
rect 198 -2320 592 1000
rect 19248 994 19744 1014
rect 19248 738 19426 994
rect 19660 738 19744 994
rect 19248 728 19744 738
rect 19402 726 19744 728
rect 30337 470 30525 471
rect 30337 466 30338 470
rect 14806 -54 15288 308
rect 22814 244 23246 286
rect 22814 200 23030 244
rect 18770 184 19414 200
rect 18770 0 19172 184
rect 19068 -36 19172 0
rect 19386 -36 19414 184
rect 22634 28 23030 200
rect 23242 28 23246 244
rect 26866 276 27258 324
rect 22634 22 23246 28
rect 26498 190 26678 200
rect 26866 190 26984 276
rect 22634 0 22814 22
rect 26498 20 26984 190
rect 27214 20 27258 276
rect 26498 0 27258 20
rect 26544 -16 27258 0
rect 19068 -46 19414 -36
rect 26866 -40 27258 -16
rect 30276 256 30338 466
rect 30524 466 30525 470
rect 30524 256 30700 466
rect 30276 -38 30700 256
rect 14806 -320 14912 -54
rect 14911 -336 14912 -320
rect 15180 -320 15288 -54
rect 15180 -336 15181 -320
rect 14911 -337 15181 -336
rect 28046 -1636 28610 -1632
rect 28046 -1998 28208 -1636
rect 28442 -1998 28610 -1636
rect 28046 -2030 28610 -1998
rect 27940 -2320 28838 -2030
rect 22 -2464 28838 -2320
rect 22 -2952 28532 -2464
rect 198 -2986 592 -2952
use sky130_fd_pr__nfet_01v8_EA9ZG2  sky130_fd_pr__nfet_01v8_EA9ZG2_0
timestamp 1724397959
transform 0 1 23920 -1 0 181
box -221 -310 221 310
use sky130_fd_pr__nfet_01v8_EA9ZG2  sky130_fd_pr__nfet_01v8_EA9ZG2_1
timestamp 1724397959
transform 0 1 19982 -1 0 85
box -221 -310 221 310
use sky130_fd_pr__pfet_01v8_EDT3T7  sky130_fd_pr__pfet_01v8_EDT3T7_0
timestamp 1724397959
transform 0 1 27729 -1 0 175
box -221 -319 221 319
<< labels >>
flabel metal4 s 30362 0 30542 200 0 FreeSans 960 0 0 0 ua[0]
port 3 nsew signal bidirectional
flabel metal4 s 26498 0 26678 200 0 FreeSans 960 0 0 0 ua[1]
port 4 nsew signal bidirectional
flabel metal4 s 22634 0 22814 200 0 FreeSans 960 0 0 0 ua[2]
port 5 nsew signal bidirectional
flabel metal4 s 18770 0 18950 200 0 FreeSans 960 0 0 0 ua[3]
port 6 nsew signal bidirectional
flabel metal4 s 14906 0 15086 200 0 FreeSans 960 0 0 0 ua[4]
port 7 nsew signal bidirectional
flabel metal4 200 1000 600 44152 1 FreeSans 400 0 0 0 VDPWR
port 51 nsew power bidirectional
flabel metal4 800 1000 1200 44152 1 FreeSans 400 0 0 0 VGND
port 52 nsew ground bidirectional
<< properties >>
string FIXED_BBOX 0 0 32200 45152
<< end >>
