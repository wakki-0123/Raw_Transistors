magic
tech sky130A
magscale 1 2
timestamp 1724397959
<< error_p >>
rect -29 172 29 178
rect -29 138 -17 172
rect -29 132 29 138
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect -29 -178 29 -172
<< pwell >>
rect -221 -310 221 310
<< nmos >>
rect -25 -100 25 100
<< ndiff >>
rect -83 88 -25 100
rect -83 -88 -71 88
rect -37 -88 -25 88
rect -83 -100 -25 -88
rect 25 88 83 100
rect 25 -88 37 88
rect 71 -88 83 88
rect 25 -100 83 -88
<< ndiffc >>
rect -71 -88 -37 88
rect 37 -88 71 88
<< psubdiff >>
rect -185 240 -89 274
rect 89 240 185 274
rect -185 178 -151 240
rect 151 178 185 240
rect -185 -240 -151 -178
rect 151 -240 185 -178
rect -185 -274 -89 -240
rect 89 -274 185 -240
<< psubdiffcont >>
rect -89 240 89 274
rect -185 -178 -151 178
rect 151 -178 185 178
rect -89 -274 89 -240
<< poly >>
rect -33 172 33 188
rect -33 138 -17 172
rect 17 138 33 172
rect -33 122 33 138
rect -25 100 25 122
rect -25 -122 25 -100
rect -33 -138 33 -122
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -33 -188 33 -172
<< polycont >>
rect -17 138 17 172
rect -17 -172 17 -138
<< locali >>
rect -185 240 -89 274
rect 89 240 185 274
rect -185 178 -151 240
rect 151 178 185 240
rect -33 138 -17 172
rect 17 138 33 172
rect -71 88 -37 104
rect -71 -104 -37 -88
rect 37 88 71 104
rect 37 -104 71 -88
rect -33 -172 -17 -138
rect 17 -172 33 -138
rect -185 -240 -151 -178
rect 151 -240 185 -178
rect -185 -274 -89 -240
rect 89 -274 185 -240
<< viali >>
rect -17 138 17 172
rect -71 -88 -37 88
rect 37 -88 71 88
rect -17 -172 17 -138
<< metal1 >>
rect -29 172 29 178
rect -29 138 -17 172
rect 17 138 29 172
rect -29 132 29 138
rect -77 88 -31 100
rect -77 -88 -71 88
rect -37 -88 -31 88
rect -77 -100 -31 -88
rect 31 88 77 100
rect 31 -88 37 88
rect 71 -88 77 88
rect 31 -100 77 -88
rect -29 -138 29 -132
rect -29 -172 -17 -138
rect 17 -172 29 -138
rect -29 -178 29 -172
<< properties >>
string FIXED_BBOX -168 -257 168 257
string gencell sky130_fd_pr__nfet_01v8
string library sky130
string parameters w 1.0 l 0.25 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__nfet_01v8 sky130_fd_pr__nfet_01v8_lvt  sky130_fd_bs_flash__special_sonosfet_star  sky130_fd_pr__nfet_g5v0d10v5 sky130_fd_pr__nfet_05v0_nvt  sky130_fd_pr__nfet_03v3_nvt} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
