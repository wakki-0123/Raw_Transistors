* NGSPICE file created from tt_um_wakki_0123_Raw_Transistors.ext - technology: sky130A

.subckt sky130_fd_pr__nfet_01v8_EA9ZG2 a_25_n100# a_n33_n188# a_n185_n274# a_n83_n100#
X0 a_25_n100# a_n33_n188# a_n83_n100# a_n185_n274# sky130_fd_pr__nfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.25
.ends

.subckt sky130_fd_pr__pfet_01v8_EDT3T7 a_25_n100# w_n221_n319# a_n83_n100# a_n33_n197#
X0 a_25_n100# a_n33_n197# a_n83_n100# w_n221_n319# sky130_fd_pr__pfet_01v8 ad=0.29 pd=2.58 as=0.29 ps=2.58 w=1 l=0.25
.ends

.subckt tt_um_wakki_0123_Raw_Transistors clk ena rst_n ua[0] ua[1] ua[2] ua[3] ua[4]
+ ua[5] ua[6] ua[7] ui_in[0] ui_in[1] ui_in[2] ui_in[3] ui_in[4] ui_in[5] ui_in[6]
+ ui_in[7] uio_in[0] uio_in[1] uio_in[2] uio_in[3] uio_in[4] uio_in[5] uio_in[6] uio_in[7]
+ uio_oe[0] uio_oe[1] uio_oe[2] uio_oe[3] uio_oe[4] uio_oe[5] uio_oe[6] uio_oe[7]
+ uio_out[0] uio_out[1] uio_out[2] uio_out[3] uio_out[4] uio_out[5] uio_out[6] uio_out[7]
+ uo_out[0] uo_out[1] uo_out[2] uo_out[3] uo_out[4] uo_out[5] uo_out[6] uo_out[7]
+ VDPWR VGND
Xsky130_fd_pr__nfet_01v8_EA9ZG2_0 ua[4] ua[2] VGND ua[0] sky130_fd_pr__nfet_01v8_EA9ZG2
Xsky130_fd_pr__nfet_01v8_EA9ZG2_1 ua[4] ua[3] VGND ua[0] sky130_fd_pr__nfet_01v8_EA9ZG2
Xsky130_fd_pr__pfet_01v8_EDT3T7_0 ua[4] VDPWR ua[0] ua[1] sky130_fd_pr__pfet_01v8_EDT3T7
.ends

