magic
tech sky130A
magscale 1 2
timestamp 1724397959
<< error_p >>
rect -29 181 29 187
rect -29 147 -17 181
rect -29 141 29 147
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect -29 -187 29 -181
<< nwell >>
rect -221 -319 221 319
<< pmos >>
rect -25 -100 25 100
<< pdiff >>
rect -83 88 -25 100
rect -83 -88 -71 88
rect -37 -88 -25 88
rect -83 -100 -25 -88
rect 25 88 83 100
rect 25 -88 37 88
rect 71 -88 83 88
rect 25 -100 83 -88
<< pdiffc >>
rect -71 -88 -37 88
rect 37 -88 71 88
<< nsubdiff >>
rect -185 249 -89 283
rect 89 249 185 283
rect -185 187 -151 249
rect 151 187 185 249
rect -185 -249 -151 -187
rect 151 -249 185 -187
rect -185 -283 -89 -249
rect 89 -283 185 -249
<< nsubdiffcont >>
rect -89 249 89 283
rect -185 -187 -151 187
rect 151 -187 185 187
rect -89 -283 89 -249
<< poly >>
rect -33 181 33 197
rect -33 147 -17 181
rect 17 147 33 181
rect -33 131 33 147
rect -25 100 25 131
rect -25 -131 25 -100
rect -33 -147 33 -131
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -33 -197 33 -181
<< polycont >>
rect -17 147 17 181
rect -17 -181 17 -147
<< locali >>
rect -185 249 -89 283
rect 89 249 185 283
rect -185 187 -151 249
rect 151 187 185 249
rect -33 147 -17 181
rect 17 147 33 181
rect -71 88 -37 104
rect -71 -104 -37 -88
rect 37 88 71 104
rect 37 -104 71 -88
rect -33 -181 -17 -147
rect 17 -181 33 -147
rect -185 -249 -151 -187
rect 151 -249 185 -187
rect -185 -283 -89 -249
rect 89 -283 185 -249
<< viali >>
rect -17 147 17 181
rect -71 -88 -37 88
rect 37 -88 71 88
rect -17 -181 17 -147
<< metal1 >>
rect -29 181 29 187
rect -29 147 -17 181
rect 17 147 29 181
rect -29 141 29 147
rect -77 88 -31 100
rect -77 -88 -71 88
rect -37 -88 -31 88
rect -77 -100 -31 -88
rect 31 88 77 100
rect 31 -88 37 88
rect 71 -88 77 88
rect 31 -100 77 -88
rect -29 -147 29 -141
rect -29 -181 -17 -147
rect 17 -181 29 -147
rect -29 -187 29 -181
<< properties >>
string FIXED_BBOX -168 -266 168 266
string gencell sky130_fd_pr__pfet_01v8
string library sky130
string parameters w 1.0 l 0.25 m 1 nf 1 diffcov 100 polycov 100 guard 1 glc 1 grc 1 gtc 1 gbc 1 tbcov 100 rlcov 100 topc 1 botc 1 poverlap 0 doverlap 1 lmin 0.15 wmin 0.42 compatible {sky130_fd_pr__pfet_01v8  sky130_fd_pr__pfet_01v8_lvt sky130_fd_pr__pfet_01v8_hvt  sky130_fd_pr__pfet_g5v0d10v5} full_metal 1 viasrc 100 viadrn 100 viagate 100 viagb 0 viagr 0 viagl 0 viagt 0
<< end >>
