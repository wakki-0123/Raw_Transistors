VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO tt_um_wakki-0123_Raw_Transistors
  CLASS BLOCK ;
  FOREIGN tt_um_wakki-0123_Raw_Transistors ;
  ORIGIN 0.000 0.000 ;
  SIZE 161.000 BY 225.760 ;
  PIN ua[0]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 151.810 0.000 152.710 1.000 ;
    END
  END ua[0]
  PIN ua[1]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.250000 ;
    PORT
      LAYER met4 ;
        RECT 132.490 0.000 133.390 1.000 ;
    END
  END ua[1]
  PIN ua[2]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.250000 ;
    PORT
      LAYER met4 ;
        RECT 113.170 0.000 114.070 1.000 ;
    END
  END ua[2]
  PIN ua[3]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.250000 ;
    PORT
      LAYER met4 ;
        RECT 93.850 0.000 94.750 1.000 ;
    END
  END ua[3]
  PIN ua[4]
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 0.870000 ;
    PORT
      LAYER met4 ;
        RECT 74.530 0.000 75.430 1.000 ;
    END
  END ua[4]
  PIN VDPWR
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER met4 ;
        RECT 1.000 5.000 3.000 220.760 ;
    END
  END VDPWR
  PIN VGND
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER met4 ;
        RECT 4.000 5.000 6.000 220.760 ;
    END
  END VGND
  OBS
      LAYER pwell ;
        RECT 98.360 -0.680 101.460 1.530 ;
        RECT 118.050 -0.200 121.150 2.010 ;
      LAYER nwell ;
        RECT 137.050 -0.230 140.240 1.980 ;
      LAYER li1 ;
        RECT 74.560 0.000 152.620 4.970 ;
        RECT 95.860 -0.180 96.930 0.000 ;
        RECT 74.560 -1.680 75.900 -0.270 ;
        RECT 98.540 -0.330 98.710 0.000 ;
        RECT 101.110 -0.330 101.280 0.000 ;
        RECT 118.230 -0.020 120.970 0.000 ;
        RECT 137.230 -0.050 140.060 0.000 ;
        RECT 98.540 -0.500 101.280 -0.330 ;
        RECT 141.040 -9.990 142.210 -8.180 ;
      LAYER met1 ;
        RECT 74.510 0.000 153.770 5.030 ;
        RECT 95.810 -0.180 96.980 0.000 ;
        RECT 74.530 -0.270 75.930 -0.210 ;
        RECT 95.830 -0.240 96.960 -0.180 ;
        RECT 99.490 -0.270 100.390 0.000 ;
        RECT 118.190 -0.110 121.060 0.000 ;
        RECT 137.200 -0.110 140.070 0.000 ;
        RECT 74.510 -1.130 75.950 -0.270 ;
        RECT 98.520 -0.570 101.390 -0.270 ;
        RECT 74.510 -1.680 76.000 -1.130 ;
        RECT 74.530 -1.740 76.000 -1.680 ;
        RECT 74.570 -1.880 76.000 -1.740 ;
        RECT 99.270 -1.880 100.540 -0.570 ;
        RECT 74.570 -1.960 100.540 -1.880 ;
        RECT 118.950 -1.960 120.430 -0.110 ;
        RECT 74.570 -2.020 120.430 -1.960 ;
        RECT 138.020 -2.020 139.470 -0.110 ;
        RECT 74.570 -2.660 139.470 -2.020 ;
        RECT 74.570 -2.810 100.540 -2.660 ;
        RECT 118.930 -2.700 139.470 -2.660 ;
        RECT 138.020 -2.750 139.470 -2.700 ;
        RECT 74.570 -2.830 76.000 -2.810 ;
        RECT 99.270 -2.840 100.540 -2.810 ;
        RECT 141.180 -3.710 142.260 0.000 ;
        RECT 141.110 -5.430 142.260 -3.710 ;
        RECT 141.110 -8.120 142.240 -5.430 ;
        RECT 141.010 -8.180 142.240 -8.120 ;
        RECT 140.990 -9.990 142.260 -8.180 ;
        RECT 141.010 -10.050 142.240 -9.990 ;
      LAYER met2 ;
        RECT 74.560 0.000 152.620 5.020 ;
        RECT 74.560 -1.730 75.900 -0.220 ;
        RECT 95.860 -0.230 96.930 0.000 ;
        RECT 141.040 -10.040 142.210 -8.130 ;
      LAYER met3 ;
        RECT 74.510 0.000 152.670 4.995 ;
        RECT 95.810 -0.205 96.980 0.000 ;
        RECT 74.510 -1.705 75.950 -0.245 ;
        RECT 140.990 -10.015 142.260 -8.155 ;
      LAYER met4 ;
        RECT 0.110 4.600 0.600 10.220 ;
        RECT 0.990 4.600 2.960 5.000 ;
        RECT 3.400 4.600 3.600 10.220 ;
        RECT 6.400 4.600 153.500 10.220 ;
        RECT 0.110 1.400 153.500 4.600 ;
        RECT 0.110 0.000 74.130 1.400 ;
        RECT 75.830 0.000 93.450 1.400 ;
        RECT 95.150 0.000 112.770 1.400 ;
        RECT 114.470 0.000 132.090 1.400 ;
        RECT 133.790 0.000 151.410 1.400 ;
        RECT 153.110 0.000 153.500 1.400 ;
        RECT 0.990 -11.600 2.960 0.000 ;
        RECT 74.030 -1.600 76.440 0.000 ;
        RECT 95.340 -0.230 97.070 0.000 ;
        RECT 132.720 -0.080 136.290 0.000 ;
        RECT 134.330 -0.200 136.290 -0.080 ;
        RECT 151.380 -0.190 153.500 0.000 ;
        RECT 74.555 -1.685 75.905 -1.600 ;
        RECT 140.230 -10.150 143.050 -8.160 ;
        RECT 139.700 -11.600 144.190 -10.150 ;
        RECT 0.110 -12.320 144.190 -11.600 ;
        RECT 0.110 -14.760 142.660 -12.320 ;
        RECT 0.990 -14.930 2.960 -14.760 ;
  END
END tt_um_wakki-0123_Raw_Transistors
END LIBRARY

